magic
tech sky130A
magscale 1 2
timestamp 1729233363
<< viali >>
rect 2764 3991 2798 4045
rect 2867 2788 2903 2857
rect 1594 2347 1628 2389
rect 3713 1278 3764 1312
<< metal1 >>
rect 2758 4045 3776 4057
rect 2758 3991 2764 4045
rect 2798 3991 3776 4045
rect 2758 3966 3776 3991
rect 3434 3754 3444 3828
rect 3510 3754 3520 3828
rect 2664 3396 3001 3430
rect 3444 3386 3509 3754
rect 2861 2864 2909 2869
rect 1586 2857 2910 2864
rect 1586 2788 2867 2857
rect 2903 2788 2910 2857
rect 1586 2776 2910 2788
rect 1587 2389 1634 2776
rect 1587 2347 1594 2389
rect 1628 2347 1634 2389
rect 1694 2566 2773 2679
rect 1694 2367 1728 2566
rect 1587 2335 1634 2347
rect 2367 1670 2377 1722
rect 2429 1670 2439 1722
rect 2712 1401 2771 2566
rect 3213 1401 3247 1641
rect 2712 1369 3247 1401
rect 3701 1312 3776 3966
rect 3701 1278 3713 1312
rect 3764 1278 3776 1312
rect 3701 1272 3776 1278
rect 2594 1191 2846 1237
rect 2594 470 2661 1191
rect 2782 542 2792 594
rect 2844 542 2854 594
rect 2375 423 2661 470
rect 2594 422 2661 423
<< via1 >>
rect 3444 3754 3510 3828
rect 2377 1670 2429 1722
rect 2792 542 2844 594
<< metal2 >>
rect 2567 3828 3510 3850
rect 2567 3754 3444 3828
rect 2567 3753 3510 3754
rect 3444 3744 3510 3753
rect 2377 1722 2429 1732
rect 2429 1670 2652 1722
rect 2377 1660 2429 1670
rect 2590 594 2652 1670
rect 2792 594 2844 604
rect 2590 542 2792 594
rect 2792 532 2844 542
use nmos  nmos_0
timestamp 1729173821
transform 1 0 2990 0 1 628
box -290 -704 978 690
use nmosout  nmosout_0
timestamp 1729222233
transform 1 0 1692 0 -1 3756
box -176 -507 1106 460
use pmoscs  pmoscs_0
timestamp 1729153036
transform 1 0 1736 0 1 458
box -178 -820 820 2052
use pmosout  pmosout_0
timestamp 1729186532
transform 1 0 3007 0 1 3029
box -176 -1590 622 574
<< end >>
