magic
tech sky130A
magscale 1 2
timestamp 1729186532
<< nwell >>
rect -176 -1590 622 574
<< nsubdiff >>
rect -140 440 -80 474
rect 526 440 586 474
rect -140 414 -106 440
rect 552 414 586 440
rect -140 -1520 -106 -1494
rect 552 -1520 586 -1494
rect -140 -1554 -80 -1520
rect 526 -1554 586 -1520
<< nsubdiffcont >>
rect -80 440 526 474
rect -140 -1494 -106 414
rect 552 -1494 586 414
rect -80 -1554 526 -1520
<< poly >>
rect -56 401 36 412
rect -56 367 -40 401
rect -6 367 36 401
rect -56 356 36 367
rect 6 330 36 356
rect 410 402 502 413
rect 410 368 452 402
rect 486 368 502 402
rect 410 357 502 368
rect 410 337 440 357
rect 94 -19 194 84
rect 94 -50 353 -19
rect -56 -110 36 -99
rect -56 -144 -40 -110
rect -6 -144 36 -110
rect 252 -143 352 -50
rect 410 -109 502 -98
rect 410 -143 452 -109
rect 486 -143 502 -109
rect -56 -155 36 -144
rect 6 -181 36 -155
rect 410 -154 502 -143
rect 410 -176 440 -154
rect -56 -606 36 -595
rect 94 -603 194 -486
rect 252 -599 351 -487
rect 410 -593 502 -582
rect -56 -640 -40 -606
rect -6 -640 36 -606
rect -56 -651 36 -640
rect 6 -677 36 -651
rect 410 -627 452 -593
rect 486 -627 502 -593
rect 410 -638 502 -627
rect 410 -664 440 -638
rect 252 -1027 352 -959
rect 94 -1057 352 -1027
rect 130 -1058 352 -1057
rect -56 -1120 36 -1109
rect 130 -1111 194 -1058
rect -56 -1154 -40 -1120
rect -6 -1154 36 -1120
rect -56 -1165 36 -1154
rect 6 -1191 36 -1165
rect 410 -1116 502 -1105
rect 410 -1150 452 -1116
rect 486 -1150 502 -1116
rect 410 -1161 502 -1150
rect 410 -1187 440 -1161
<< polycont >>
rect -40 367 -6 401
rect 452 368 486 402
rect -40 -144 -6 -110
rect 452 -143 486 -109
rect -40 -640 -6 -606
rect 452 -627 486 -593
rect -40 -1154 -6 -1120
rect 452 -1150 486 -1116
<< locali >>
rect -140 440 -80 474
rect 526 440 586 474
rect -140 414 -106 440
rect 552 414 586 440
rect -56 367 -40 401
rect -6 367 10 401
rect 436 368 452 402
rect 486 368 502 402
rect -56 -144 -40 -110
rect -6 -144 10 -110
rect 436 -143 452 -109
rect 486 -143 502 -109
rect -56 -640 -40 -606
rect -6 -640 10 -606
rect 436 -627 452 -593
rect 486 -627 502 -593
rect -56 -1154 -40 -1120
rect -6 -1154 10 -1120
rect 436 -1150 452 -1116
rect 486 -1150 502 -1116
rect -140 -1520 -106 -1494
rect 552 -1520 586 -1494
rect -140 -1554 -80 -1520
rect 526 -1554 586 -1520
<< viali >>
rect 208 440 242 474
rect -40 367 -6 401
rect 452 368 486 402
rect -40 -144 -6 -110
rect 452 -143 486 -109
rect -40 -640 -6 -606
rect 452 -627 486 -593
rect -40 -1154 -6 -1120
rect 452 -1150 486 -1116
<< metal1 >>
rect 193 474 260 487
rect 193 440 208 474
rect 242 440 260 474
rect 193 434 260 440
rect -52 401 6 407
rect -52 367 -40 401
rect -6 367 6 401
rect 440 402 498 408
rect -52 356 6 367
rect -40 308 -6 356
rect 109 339 176 389
rect 270 339 337 389
rect 440 368 452 402
rect 486 368 498 402
rect 440 357 498 368
rect 452 308 486 357
rect -40 243 82 308
rect -62 187 -52 243
rect 4 187 82 243
rect -40 132 82 187
rect 100 81 174 83
rect 100 31 176 81
rect 100 29 174 31
rect -63 -70 -53 -14
rect 3 -70 13 -14
rect -41 -104 -7 -70
rect 100 -101 174 -100
rect -52 -110 6 -104
rect -52 -144 -40 -110
rect -6 -144 6 -110
rect -52 -155 6 -144
rect 100 -153 114 -101
rect 166 -153 176 -101
rect 100 -154 174 -153
rect -41 -194 -6 -155
rect -40 -379 82 -203
rect -52 -606 6 -600
rect -52 -640 -40 -606
rect -6 -640 6 -606
rect -52 -651 6 -640
rect -40 -695 -6 -651
rect 42 -699 71 -379
rect 100 -430 174 -428
rect 100 -480 176 -430
rect 100 -482 174 -480
rect 100 -598 174 -596
rect 100 -648 176 -598
rect 100 -650 174 -648
rect -40 -861 82 -699
rect -41 -875 82 -861
rect -41 -939 -6 -875
rect 100 -925 174 -924
rect -62 -995 -52 -939
rect 4 -995 14 -939
rect 100 -977 115 -925
rect 167 -977 177 -925
rect 100 -978 174 -977
rect 100 -1113 177 -1108
rect -52 -1120 6 -1114
rect -52 -1154 -40 -1120
rect -6 -1154 6 -1120
rect -52 -1165 6 -1154
rect -40 -1208 -6 -1165
rect 99 -1167 177 -1113
rect -40 -1274 82 -1213
rect -62 -1330 -52 -1274
rect 4 -1330 82 -1274
rect -40 -1389 82 -1330
rect 206 -1381 240 300
rect 364 132 486 308
rect 272 82 346 83
rect 271 81 281 82
rect 270 31 281 81
rect 271 30 281 31
rect 333 30 346 82
rect 452 79 486 132
rect 272 29 346 30
rect 431 23 441 79
rect 497 23 507 79
rect 268 -156 346 -97
rect 440 -109 498 -103
rect 440 -143 452 -109
rect 486 -143 498 -109
rect 440 -154 498 -143
rect 452 -203 486 -154
rect 364 -238 486 -203
rect 364 -294 446 -238
rect 502 -294 512 -238
rect 364 -379 486 -294
rect 268 -484 346 -425
rect 268 -652 346 -593
rect 374 -699 403 -379
rect 440 -593 498 -587
rect 440 -627 452 -593
rect 486 -627 498 -593
rect 440 -638 498 -627
rect 452 -699 486 -638
rect 364 -758 486 -699
rect 364 -814 443 -758
rect 499 -814 509 -758
rect 364 -875 486 -814
rect 268 -980 346 -921
rect 427 -1070 437 -1014
rect 493 -1070 503 -1014
rect 450 -1110 486 -1070
rect 272 -1111 346 -1110
rect 272 -1112 282 -1111
rect 270 -1162 282 -1112
rect 272 -1163 282 -1162
rect 334 -1163 346 -1111
rect 440 -1116 498 -1110
rect 440 -1150 452 -1116
rect 486 -1150 498 -1116
rect 440 -1161 498 -1150
rect 272 -1164 346 -1163
rect 452 -1212 486 -1161
rect 364 -1389 486 -1213
rect 109 -1470 176 -1420
rect 269 -1470 336 -1420
<< via1 >>
rect -52 187 4 243
rect -53 -70 3 -14
rect 114 -153 166 -101
rect -52 -995 4 -939
rect 115 -977 167 -925
rect -52 -1330 4 -1274
rect 281 30 333 82
rect 441 23 497 79
rect 446 -294 502 -238
rect 443 -814 499 -758
rect 437 -1070 493 -1014
rect 282 -1163 334 -1111
<< metal2 >>
rect -52 243 4 253
rect -52 177 4 187
rect 281 82 333 92
rect 281 20 333 30
rect 441 79 497 89
rect -53 -14 3 -4
rect 281 -18 332 20
rect 441 13 497 23
rect -53 -80 3 -70
rect 114 -55 332 -18
rect 114 -60 331 -55
rect 114 -101 166 -60
rect 114 -163 166 -153
rect 446 -238 502 -228
rect 446 -304 502 -294
rect 443 -758 499 -748
rect 443 -824 499 -814
rect 115 -925 167 -915
rect -52 -939 4 -929
rect -52 -1005 4 -995
rect 115 -979 167 -977
rect 115 -1027 168 -979
rect 437 -1014 493 -1004
rect 115 -1062 335 -1027
rect 283 -1101 335 -1062
rect 437 -1080 493 -1070
rect 282 -1111 335 -1101
rect 282 -1173 334 -1163
rect -52 -1274 4 -1264
rect -52 -1340 4 -1330
<< via2 >>
rect -52 187 4 243
rect 441 23 497 79
rect -53 -70 3 -14
rect 446 -294 502 -238
rect 443 -814 499 -758
rect -52 -995 4 -939
rect 437 -1070 493 -1014
rect -52 -1330 4 -1274
<< metal3 >>
rect -77 249 24 262
rect -77 171 -59 249
rect 13 171 24 249
rect -77 155 24 171
rect 431 79 507 84
rect 431 23 441 79
rect 497 23 507 79
rect 431 -9 507 23
rect -63 -14 507 -9
rect -63 -70 -53 -14
rect 3 -70 507 -14
rect -63 -78 507 -70
rect 425 -234 530 -215
rect 425 -300 442 -234
rect 515 -300 530 -234
rect 425 -322 530 -300
rect 422 -751 526 -743
rect 422 -821 436 -751
rect 514 -821 526 -751
rect 422 -841 526 -821
rect -62 -935 14 -934
rect -62 -939 15 -935
rect -62 -995 -52 -939
rect 4 -995 15 -939
rect -62 -1009 15 -995
rect -62 -1014 503 -1009
rect -62 -1070 437 -1014
rect 493 -1070 503 -1014
rect -62 -1076 503 -1070
rect -76 -1268 33 -1256
rect -76 -1336 -55 -1268
rect 14 -1336 33 -1268
rect -76 -1357 33 -1336
<< via3 >>
rect -59 243 13 249
rect -59 187 -52 243
rect -52 187 4 243
rect 4 187 13 243
rect -59 171 13 187
rect 442 -238 515 -234
rect 442 -294 446 -238
rect 446 -294 502 -238
rect 502 -294 515 -238
rect 442 -300 515 -294
rect 436 -758 514 -751
rect 436 -814 443 -758
rect 443 -814 499 -758
rect 499 -814 514 -758
rect 436 -821 514 -814
rect -55 -1274 14 -1268
rect -55 -1330 -52 -1274
rect -52 -1330 4 -1274
rect 4 -1330 14 -1274
rect -55 -1336 14 -1330
<< metal4 >>
rect -72 249 27 255
rect -72 171 -59 249
rect 13 171 27 249
rect -72 82 27 171
rect -72 81 522 82
rect -72 34 530 81
rect -70 -32 530 34
rect 428 -213 530 -32
rect 421 -234 537 -213
rect 421 -300 442 -234
rect 515 -300 537 -234
rect 421 -328 537 -300
rect 412 -751 533 -727
rect 412 -821 436 -751
rect 514 -821 533 -751
rect 412 -852 533 -821
rect 413 -1014 519 -852
rect -70 -1024 519 -1014
rect -82 -1100 519 -1024
rect -82 -1250 46 -1100
rect 413 -1102 519 -1100
rect -83 -1268 46 -1250
rect -83 -1336 -55 -1268
rect 14 -1336 46 -1268
rect -83 -1372 46 -1336
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_0
timestamp 1729178293
transform 1 0 21 0 1 220
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_1
timestamp 1729178293
transform 1 0 425 0 1 220
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_2
timestamp 1729178293
transform 1 0 21 0 1 -291
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_3
timestamp 1729178293
transform 1 0 425 0 1 -291
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_4
timestamp 1729178293
transform 1 0 21 0 1 -1301
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_5
timestamp 1729178293
transform 1 0 425 0 1 -1301
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_6
timestamp 1729178293
transform 1 0 21 0 1 -787
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_7
timestamp 1729178293
transform 1 0 425 0 1 -787
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_VQXX6L  sky130_fd_pr__pfet_01v8_VQXX6L_0
timestamp 1729179451
transform 1 0 223 0 1 -1301
box -223 -200 223 200
use sky130_fd_pr__pfet_01v8_VQXX6L  sky130_fd_pr__pfet_01v8_VQXX6L_1
timestamp 1729179451
transform 1 0 223 0 1 -787
box -223 -200 223 200
use sky130_fd_pr__pfet_01v8_VQXX6L  sky130_fd_pr__pfet_01v8_VQXX6L_2
timestamp 1729179451
transform 1 0 223 0 1 -291
box -223 -200 223 200
use sky130_fd_pr__pfet_01v8_VQXX6L  sky130_fd_pr__pfet_01v8_VQXX6L_3
timestamp 1729179451
transform 1 0 223 0 1 220
box -223 -200 223 200
<< labels >>
flabel viali 219 462 219 462 0 FreeSans 800 0 0 0 vdd
port 1 nsew
flabel metal1 227 261 227 261 0 FreeSans 800 0 0 0 s
port 2 nsew
flabel metal1 124 375 124 375 0 FreeSans 800 0 0 0 vin
port 3 nsew
flabel metal1 300 378 300 378 0 FreeSans 800 0 0 0 vip
port 4 nsew
flabel via3 -43 195 -43 195 0 FreeSans 800 0 0 0 d6
port 5 nsew
flabel metal1 467 203 467 203 0 FreeSans 800 0 0 0 out
port 6 nsew
<< end >>
