magic
tech sky130A
magscale 1 2
timestamp 1729173821
<< nmos >>
rect -144 88 -114 488
rect -144 -545 -114 -145
rect 58 -545 258 -145
rect 430 -545 630 -145
rect 802 -545 832 -145
<< ndiff >>
rect -202 476 -144 488
rect -202 100 -190 476
rect -156 100 -144 476
rect -202 88 -144 100
rect -114 476 -56 488
rect -114 100 -102 476
rect -68 100 -56 476
rect -114 88 -56 100
rect -202 -157 -144 -145
rect -202 -533 -190 -157
rect -156 -533 -144 -157
rect -202 -545 -144 -533
rect -114 -157 -56 -145
rect -114 -533 -102 -157
rect -68 -533 -56 -157
rect -114 -545 -56 -533
rect 0 -157 58 -145
rect 0 -533 12 -157
rect 46 -533 58 -157
rect 0 -545 58 -533
rect 258 -157 316 -145
rect 258 -533 270 -157
rect 304 -533 316 -157
rect 258 -545 316 -533
rect 372 -157 430 -145
rect 372 -533 384 -157
rect 418 -533 430 -157
rect 372 -545 430 -533
rect 630 -157 688 -145
rect 630 -533 642 -157
rect 676 -533 688 -157
rect 630 -545 688 -533
rect 744 -157 802 -145
rect 744 -533 756 -157
rect 790 -533 802 -157
rect 744 -545 802 -533
rect 832 -157 890 -145
rect 832 -533 844 -157
rect 878 -533 890 -157
rect 832 -545 890 -533
<< ndiffc >>
rect -190 100 -156 476
rect -102 100 -68 476
rect -190 -533 -156 -157
rect -102 -533 -68 -157
rect 12 -533 46 -157
rect 270 -533 304 -157
rect 384 -533 418 -157
rect 642 -533 676 -157
rect 756 -533 790 -157
rect 844 -533 878 -157
<< psubdiff >>
rect -290 650 -230 684
rect 918 650 978 684
rect -290 624 -256 650
rect 944 624 978 650
rect -290 -664 -256 -638
rect 944 -664 978 -638
rect -290 -698 -230 -664
rect 918 -698 978 -664
<< psubdiffcont >>
rect -230 650 918 684
rect -290 -638 -256 624
rect 944 -638 978 624
rect -230 -698 918 -664
<< poly >>
rect -206 603 -114 619
rect -206 569 -190 603
rect -156 569 -114 603
rect -206 553 -114 569
rect -144 488 -114 553
rect 802 570 894 586
rect 802 536 844 570
rect 878 536 894 570
rect 802 520 894 536
rect 802 514 832 520
rect -144 62 -114 88
rect -206 -42 -114 -26
rect -206 -76 -190 -42
rect -156 -76 -114 -42
rect -206 -92 -114 -76
rect -144 -145 -114 -92
rect 58 -73 630 50
rect 58 -107 74 -73
rect 242 -107 446 -73
rect 614 -107 630 -73
rect 58 -145 258 -107
rect 430 -145 630 -107
rect 802 -58 894 -42
rect 802 -92 844 -58
rect 878 -92 894 -58
rect 802 -108 894 -92
rect 802 -145 832 -108
rect -144 -571 -114 -545
rect 58 -583 258 -545
rect 58 -617 74 -583
rect 242 -617 258 -583
rect 58 -633 258 -617
rect 430 -583 630 -545
rect 802 -571 832 -545
rect 430 -617 446 -583
rect 614 -617 630 -583
rect 430 -633 630 -617
<< polycont >>
rect -190 569 -156 603
rect 844 536 878 570
rect -190 -76 -156 -42
rect 74 -107 242 -73
rect 446 -107 614 -73
rect 844 -92 878 -58
rect 74 -617 242 -583
rect 446 -617 614 -583
<< locali >>
rect -290 650 -230 684
rect 918 650 978 684
rect -290 624 -256 650
rect 944 624 978 650
rect -206 569 -190 603
rect -156 569 -140 603
rect 828 536 844 570
rect 878 536 894 570
rect -190 476 -156 492
rect -190 84 -156 100
rect -102 476 -68 492
rect -102 84 -68 100
rect -206 -76 -190 -42
rect -156 -76 -140 -42
rect 58 -107 74 -73
rect 242 -107 258 -73
rect 430 -107 446 -73
rect 614 -107 630 -73
rect 828 -92 844 -58
rect 878 -92 894 -58
rect -190 -157 -156 -141
rect -190 -549 -156 -533
rect -102 -157 -68 -141
rect -102 -549 -68 -533
rect 12 -157 46 -141
rect 12 -549 46 -533
rect 270 -157 304 -141
rect 270 -549 304 -533
rect 384 -157 418 -141
rect 384 -549 418 -533
rect 642 -157 676 -141
rect 642 -549 676 -533
rect 756 -157 790 -141
rect 756 -549 790 -533
rect 844 -157 878 -141
rect 844 -549 878 -533
rect 58 -617 74 -583
rect 242 -617 258 -583
rect 430 -617 446 -583
rect 614 -617 630 -583
rect -290 -664 -256 -638
rect 944 -664 978 -638
rect -290 -698 -230 -664
rect 918 -698 978 -664
<< viali >>
rect 270 650 304 684
rect -190 569 -156 603
rect 844 536 878 570
rect -190 100 -156 476
rect -102 100 -68 476
rect -190 -76 -156 -42
rect 99 -107 217 -73
rect 471 -107 589 -73
rect 844 -92 878 -58
rect -190 -533 -156 -157
rect -102 -533 -68 -157
rect 12 -533 46 -157
rect 270 -533 304 -157
rect 384 -533 418 -157
rect 642 -533 676 -157
rect 756 -533 790 -157
rect 844 -533 878 -157
rect 99 -617 217 -583
rect 471 -617 589 -583
rect 384 -698 418 -664
<< metal1 >>
rect 258 684 316 690
rect 258 650 270 684
rect 304 650 316 684
rect 258 644 316 650
rect -202 603 -144 609
rect -202 569 -190 603
rect -156 569 -144 603
rect -202 563 -144 569
rect -190 488 -156 563
rect -196 476 -150 488
rect -108 476 -62 488
rect -196 100 -190 476
rect -156 100 -102 476
rect -68 475 -62 476
rect -68 100 46 475
rect -196 88 -150 100
rect -108 88 -62 100
rect 7 50 52 88
rect 7 16 99 50
rect 270 -7 304 644
rect 832 570 890 576
rect 832 536 844 570
rect 878 536 890 570
rect 832 530 890 536
rect 844 476 878 530
rect 642 118 878 476
rect 756 100 878 118
rect 352 36 362 88
rect 414 36 427 88
rect 632 32 642 88
rect 698 32 708 88
rect -202 -42 -144 -36
rect 269 -40 419 -7
rect -202 -76 -190 -42
rect -156 -76 -144 -42
rect -202 -82 -144 -76
rect 87 -73 229 -67
rect -190 -145 -156 -82
rect -20 -145 -10 -89
rect 46 -145 56 -89
rect 87 -107 99 -73
rect 217 -107 229 -73
rect 87 -113 229 -107
rect 266 -145 276 -93
rect 328 -145 338 -93
rect 384 -145 418 -40
rect 832 -58 890 -52
rect 459 -73 601 -67
rect 459 -107 471 -73
rect 589 -107 682 -73
rect 832 -92 844 -58
rect 878 -92 890 -58
rect 832 -98 890 -92
rect 459 -113 601 -107
rect -196 -157 -150 -145
rect -108 -157 -62 -145
rect -196 -533 -190 -157
rect -156 -533 -102 -157
rect -68 -175 -62 -157
rect 6 -157 52 -145
rect 6 -175 12 -157
rect -68 -533 12 -175
rect 46 -533 52 -157
rect -196 -545 -150 -533
rect -108 -545 -62 -533
rect 6 -545 52 -533
rect 264 -157 310 -145
rect 264 -533 270 -157
rect 304 -533 310 -157
rect 264 -545 310 -533
rect 378 -157 424 -145
rect 378 -533 384 -157
rect 418 -533 424 -157
rect 378 -545 424 -533
rect 636 -157 682 -107
rect 844 -145 878 -98
rect 750 -157 796 -145
rect 838 -157 884 -145
rect 636 -533 642 -157
rect 676 -533 756 -157
rect 790 -533 844 -157
rect 878 -533 884 -157
rect 636 -545 682 -533
rect 750 -545 796 -533
rect 838 -545 884 -533
rect 87 -583 229 -577
rect 87 -617 99 -583
rect 217 -617 229 -583
rect 87 -623 229 -617
rect 384 -658 418 -545
rect 459 -583 601 -577
rect 459 -617 471 -583
rect 589 -617 601 -583
rect 459 -623 601 -617
rect 372 -664 430 -658
rect 372 -698 384 -664
rect 418 -698 430 -664
rect 372 -704 430 -698
<< via1 >>
rect 362 36 414 88
rect 642 32 698 88
rect -10 -145 46 -89
rect 276 -145 328 -93
<< metal2 >>
rect 362 88 414 98
rect 362 -7 414 36
rect 642 88 698 98
rect 642 22 698 32
rect 276 -39 414 -7
rect -10 -89 46 -79
rect -10 -155 46 -145
rect 276 -93 329 -39
rect 328 -145 329 -93
rect 276 -155 328 -145
<< via2 >>
rect 642 32 698 88
rect -10 -145 46 -89
<< metal3 >>
rect 632 88 708 93
rect 632 32 642 88
rect 698 32 708 88
rect 632 7 708 32
rect -20 -55 708 7
rect -20 -89 56 -55
rect -20 -145 -10 -89
rect 46 -145 56 -89
rect -20 -150 56 -145
use sky130_fd_pr__nfet_01v8_6C7GGL  sky130_fd_pr__nfet_01v8_6C7GGL_0
timestamp 1729155829
transform 1 0 817 0 1 288
box -73 -226 73 226
use sky130_fd_pr__nfet_01v8_8UMB6F  sky130_fd_pr__nfet_01v8_8UMB6F_0
timestamp 1729158240
transform 1 0 344 0 1 288
box -344 -288 344 288
<< labels >>
flabel metal1 288 228 288 228 0 FreeSans 320 0 0 0 S3
flabel metal1 30 231 30 231 0 FreeSans 320 0 0 0 D3
flabel space 400 223 400 223 0 FreeSans 320 0 0 0 S4
flabel metal1 667 217 667 217 0 FreeSans 320 0 0 0 D4
flabel viali 287 -309 287 -309 0 FreeSans 320 0 0 0 S4
flabel viali 30 -318 30 -318 0 FreeSans 320 0 0 0 D4
flabel viali 400 -333 400 -333 0 FreeSans 320 0 0 0 S3
flabel viali 657 -337 657 -337 0 FreeSans 320 0 0 0 D3
flabel viali 399 -681 399 -681 0 FreeSans 1600 0 0 0 gnd
port 1 nsew
flabel via1 382 67 382 67 0 FreeSans 1600 0 0 0 rs
port 2 nsew
flabel metal1 29 42 29 42 0 FreeSans 1600 0 0 0 d3
port 3 nsew
flabel via2 669 54 669 54 0 FreeSans 1600 0 0 0 d4
port 4 nsew
<< end >>
