magic
tech sky130A
magscale 1 2
timestamp 1729054082
<< metal1 >>
rect 322 2354 1673 2536
rect 405 2107 447 2354
rect 826 2117 868 2354
rect 1250 2113 1292 2354
rect 509 1914 613 1920
rect 509 1859 517 1914
rect 605 1859 613 1914
rect 1494 1912 1598 1920
rect 652 1871 1019 1905
rect 1074 1872 1439 1905
rect 509 1851 613 1859
rect 1494 1858 1502 1912
rect 1591 1858 1598 1912
rect 1494 1851 1598 1858
rect 407 1438 449 1790
rect 827 1438 869 1778
rect 1248 1438 1290 1777
rect 310 1256 1661 1438
<< via1 >>
rect 517 1859 605 1914
rect 1502 1858 1591 1912
<< metal2 >>
rect 509 1914 1598 1920
rect 509 1859 517 1914
rect 605 1912 1598 1914
rect 605 1859 1502 1912
rect 509 1858 1502 1859
rect 1591 1858 1598 1912
rect 509 1852 1598 1858
use inverter  x1
timestamp 1729052800
transform 1 0 423 0 1 1306
box -53 21 369 1147
use inverter  x2
timestamp 1729052800
transform 1 0 844 0 1 1306
box -53 21 369 1147
use inverter  x3
timestamp 1729052800
transform 1 0 1265 0 1 1306
box -53 21 369 1147
<< labels >>
flabel metal1 400 2464 400 2464 0 FreeSans 800 0 0 0 VDD
port 1 nsew
flabel metal1 400 1316 400 1316 0 FreeSans 800 0 0 0 GND
port 2 nsew
flabel metal2 826 1888 826 1891 0 FreeSans 800 0 0 0 OUT
port 3 nsew
<< end >>
